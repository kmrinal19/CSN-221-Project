module memory ();
    reg [31:0] memory[0:1023];
endmodule