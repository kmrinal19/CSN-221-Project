module PC();
integer pc;
initial pc=0;
endmodule